----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 28.12.2022 22:25:33
-- Design Name: 
-- Module Name: affichage - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity affichage is
    Port ( RESET : in STD_LOGIC;
           clk : in STD_LOGIC;
           Nb1 : in STD_LOGIC_VECTOR (15 downto 0);
           Nb2 : in STD_LOGIC_VECTOR (15 downto 0);
           Resultat : in STD_LOGIC_VECTOR (15 downto 0);
           Progress : in STD_LOGIC_VECTOR (1 downto 0));
end affichage;

architecture Behavioral of affichage is

begin


end Behavioral;
